library IEEE ;
USE IEEE.std_logic_1164.all ; --std_logic_1164不要忘

entity dff1 is
	Port(CL,CK,T: in std_logic;
	     Q,Qbar: out std_logic);
		  
end dff1 ;

architecture arch of dff1 is
begin
	Process(cl,ck)
	begin
		if t='1' then 
		elsif reisng then
		if t = 1 t te p 
		ese ruell
		endi f
		q<=tmp
		